    00     �%  6          �  �%       h  �6  (   0   `           $                                                                                                                                                                                                                  ���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������uxx�^``�WWW�VVV�VVV�VVV�VVV�VVV�VVV�VVV�VVV�VVV�VVV�VVV�VVV�VVV�VVV�WWW�^``�txx�����������������������������������������������������������������������������������������������������]^^�2�H�n  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �o  �I�2�\]]���������������������������������������������������������������������������������tvv�.�u  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �� �� �� �� ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �v  �.�suu���������������������������������������������������������������������OOO�H��  �� ��  ��  ��  ��  ��  ��  ��  �� �� �� �� �� �� �� �� �� ��  ��  ��  ��  ��  ��  ��  ��  �� ��  �J�MMM�������������������������������������������������������������POO�Z  �� ��  ��  ��  ��  ��  ��  �� �� �f�5�%�)'�02�47�25�--�&�*�I�� �� ��  ��  ��  ��  ��  ��  ��  ���\  �MMM�����������������������������������������������������suu�K��  ��  ��  ��  ��  ��  �� �� �E�#�<@�^b�su�|~� ��� �� ��~ ��xz�jm�NS�+,�*�t �� ��  ��  ��  ��  ��  ��  �� �M�qss�������������������������������������������������0��  ��  ��  ��  ��  ��  ���c� �GL�su�� ��� ��� �� �� �� �� �� �� ��� ��� ��| ~�ad�-/�1�� ����  ��  ��  ��  ��  ��  �1���������������������������������������������[\\�y  ��  ��  ��  ��  ��  �� �;�.1�mo�� ��� �� �� �� �� �� �� �� �� �� �� �� �� ��� ��|~�PS� � ����  ��  ��  ��  ��  �|  �YYY�����������������������������������������3��  ��  ��  ��  ��  �� �0�>B�z|�� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��� ��dg�!�s �� ��  ��  ��  ��  ��  �3�����������������������������������������L��  ��  ��  ��  �� �5�AD�}�� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��� ��il� �� �� ��  ��  ��  ��  �N�������������������������������������qtt�u  ��  ��  ��  ���S�48�|}�� �� �� �� ��~ ��} �~ �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��� ��ad� �� ��  ��  ��  ��  �y  �nqq���������������������������������Z[[��  ��  ��  �� �� �"�st�� �� �� �� ������`�������M�� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��� ��IM�:�� ��  ��  ��  ��  �XXX���������������������������������SRR��  ��  ��  �� �2�UY�� �� �� �� �� ���
����������˚�� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��� ��y{�''�� �� ��  ��  ��  �POO���������������������������������RQQ��  ��  ��  �� �('�z|� �� �� �� �� ���
����������˙��~ �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��� ��WZ�5�� ��  ��  ��  �ONN���������������������������������RQQ��  ��  ���B�OS�� �� �� �� �� �� ���
����������˙��~ �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��� ��xz�$ �� ��  ��  ��  �PNN���������������������������������RQQ��  ��  �� �$�or�� �� �� �� �� �� ���
����������˙��~ �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��� ��>C�b ��  ��  ��  �ONN���������������������������������RQQ��  ��  �� �**�}~� �� �� �� �� �� ���
����������˙��~ �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��� ��[`�7����  ��  �ONN���������������������������������RQQ��  ��  �n �;@�� �� �� �� �� �� �� ���
����������ʙ��} �~ ��~ ��~ ��~ ��~ �� �� �� �� �� �� �� �� �� �� �� ��� ��mq�'�� ��  ��  �ONN���������������������������������RQQ��  ��  �V�IO�� �� �� �� �� �� �� ���
����������Ҩ���$���$���$���$���$��� ��������} � �� �� �� �� �� �� �� ��� ��vx�$�� ��  ��  �ONN���������������������������������RQQ��  ��  �J�QV�� �� �� �� �� �� �� ���
������������������������������������������Ϣ���P���	��~ �� �� �� �� �� �� �� ��y |�% �� ��  ��  �ONN���������������������������������RQQ��  ��  �J�QV�� �� �� �� �� �� �� ���
��������������������������������������������������Ì���
�� �� �� �� �� �� �� ��y |�% �� ��  ��  �ONN���������������������������������RQQ��  ��  �T�JO�� �� �� �� �� �� �� ���
����������Ԭ���/���0���0���0���1���>���j���������������c��~ � �� �� �� �� ��� ��wy�%�� ��  ��  �ONN���������������������������������RQQ��  ��  �k �=A�� �� �� �� �� �� �� ���
����������ʙ��} �~ ��~ ��~ ��} ��} �} ~��!����������������� �� �� �� �� ��� ��nq�'�� ��  ��  �ONN���������������������������������RQQ��  ��  �� �+,�}� �� �� �� �� �� ���
����������˙��~ �� �� �� �� �� �� ��} ~��v�����������+��~ �� �� �� �� ��� ��]a�5�� ��  ��  �ONN���������������������������������RQQ��  ��  �� �$�qs�� �� �� �� �� �� ���
����������˙��~ �� �� �� �� �� �� ��} ��^�����������8��} � �� �� �� ��� ��AE�^ ��  ��  ��  �ONN���������������������������������RQQ��  ��  �� �>�RV�� �� �� �� �� �� ���
����������˙��~ �� �� �� �� �� �� ��} �������������+��~ �� �� �� �� ��y{�&"�� ��  ��  ��  �ONN���������������������������������RQQ��  ��  ��  �� �**�|}� �� �� �� �� ���
����������ʙ��| ~�} ~�} ~�} ~�} �} �} ��1����������޿����� �� �� �� ��� ��Z^�1�� ��  ��  ��  �ONN���������������������������������SRR��  ��  ��  �� �.�Y\�� �� �� �� �� ���
����������ݽ���Z���[���[���[���\���c�������������������]��~ � �� �� �� ��{|�**�� �� ��  ��  ��  �POO���������������������������������YZZ��  ��  ��  �� �� �$"�uw�� �� �� �� ���
���������������������������������������������������{����� �� �� �� ��� ��NR�5����  ��  ��  ��  �VVV���������������������������������nqq�x  ��  ��  ��  �� �J�9=�}� �� �� �����ȓ������������������������������ܻ��Ӫ�������8����� �� �� �� ��� ��gi� �� �� ��  ��  ��  �{  �knn�������������������������������������P��  ��  ��  ��  �� �/�GK�~ �� �� �� ������������������������
��������} �~ �� �� �� �� ��� ��np�" �y ����  ��  ��  �� �R�����������������������������������������4��  ��  ��  ��  �� �� �)�FJ�}~�� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��� ��jl�$"�g �� ��  ��  ��  ��  ��  �3�����������������������������������������UUU��  ��  ��  ��  ��  �� �� �3�58�rt�� ��� �� �� �� �� �� �� �� �� �� �� �� �� ��� ��~��X[� �r �� ��  ��  ��  ��  �� ��  �SRR���������������������������������������������2��  ��  ��  ��  ��  �� ���V�"�PT�wy�� ��� ��� �� �� �� �� �� �� ��� ��� ��~ ��hj�47�*	�� ����  ��  ��  ��  ��  ��  �2�������������������������������������������������ikk�R  �� ��  ��  ��  ��  ��  ���� �;�$ �CH�eh�wy�~ ��� ��� ��� �� ��{ }�or�UY�13�%�g�� �� ��  ��  ��  ��  ��  ��  �T  �fih�����������������������������������������������������FDE�e  �� ��  ��  ��  ��  ��  ��  �� �� �V�+�$�,-�48�9>�8<�03�'%�$�;�z �� �� ��  ��  ��  ��  ��  ��  ��  �h  �EBB�������������������������������������������������������������FDD�T  ��  �� ��  ��  ��  ��  ��  ��  ��  �� �� �� �| �r �u �� �� �� ��  ��  ��  ��  ��  ��  ��  ��  �� ��  �V  �DBB���������������������������������������������������������������������hjj�1��  ��  �� �� ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �� ��  ��  �2�ghh���������������������������������������������������������������������������������PPP�2�S�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �T�2�OOO�����������������������������������������������������������������������������������������������������ehh�RQQ�KHH�JGG�JGG�JGG�JGG�JGG�JGG�JGG�JGG�JGG�JGG�JGG�JGG�JGG�JGG�KHH�RPP�egg������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=                                                                                                                                                                                                ������  ������                                                                                                                                                                                                                                                                                                                                                                  ������  ������  (       @                             ssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssss����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������lLL�l!!�w�z�z�{�|�|�|�{�{�z�z�w�m!!�lLL���������������������������������������������������������eFF����  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ���eEE���������������������������������������������`--��  ��  ��  ��  ��  �� ���_�N �I(�J&�R�k����  ��  ��  ��  ��  ��  �`,,�������������������������������������fFF��  ��  ��  ��  �� �q�D-�UX�lq�w |�z �z ~�t y�ek�MK�I����  ��  ��  ��  ��  �fEE������������������������������������  ��  ��  �� �H�X\�{ ~�� ��� �� �� �� �� ��� ��� ��sx�IH�`�� ��  ��  ��  �������������������������������lJJ��  ��  ��  �� �A'�lq�� �� �� �� �� �� �� �� �� �� ��� �� ��Y]�T�� ��  ��  ��  �kHH�������������������������o  ��  ��  �� �E �nr�� �� ������ �� �� �� �� �� �� �� �� ��� ��W[�d�� ��  ��  �p�������������������������{��  ��  �d�^b�� �� ��~ ���Y��ʙ�����~ �� �� �� �� �� �� �� �� �� ��GC����  ��  �|�������������������������~��  �� �D8�~ �� �� ��~ �Ċ�������*��~ �� �� �� �� �� �� �� �� ��� ��ot�N�� ��  ��������������������������~��  �r	�_d�� �� �� ��~ �Ċ�������*��~ �� �� �� �� �� �� �� �� �� ��� ��HB�� ��  ����������������������������  �N�u y� �� �� ��~ �Ċ�������*��~ �� �� �� �� �� �� �� �� �� ��� ��]b�{��  �����������������������������  �F0�} �� �� �� ��~ �Ċ�������,�� ����������} �~ �� �� �� �� ��� ��mr�]��  ������������������������������  �G;� �� �� �� ��~ �É������ܻ��խ��֮��խ��͛���e�����~ �� �� �� ��� ��s x�S��  ������������������������������  �G;�� �� �� �� ��~ �É����������ڷ��۸��ܻ����������ۺ�����~ �� �� ��� ��s y�R��  ������������������������������  �F1�~ �� �� �� ��~ �Ċ�������/���������������x�������z��~ �� �� ��� ��ms�]��  �����������������������������  �M�uz� �� �� ��~ �Ċ�������*��~ �� �� ��~ ���������ٴ����� �� ��� ��^c�x��  ��������������������������~��  �p
�`e�� �� �� ��~ �Ċ�������*��} �~ ��~ ��} ��������ٴ����� �� ��� ��IC�� ��  ��������������������������~��  �� �E:�~ �� �� ��~ �ĉ�������9�����������������������x��~ �� ��� ��qv�M�� ��  ��������������������������{��  ��  �`�`e�� �� ��~ ��É������������������������������ְ�����~ �� �� ��HF����  ��  �|�������������������������p��  ��  �� �C#�pu�� ��~ ���I��Č��Č��Ō��Ō��Ê���|���P�����~ �� ��� ��[_�_�� ��  ��  �p�������������������������kGG��  ��  ��  ���A,�ot�� ��~ ��~ ��~ ��~ ��~ ��} �} �} �~ ��� ��� ��]a�P�� ��  ��  ��  �jEE��������������������������������  ��  ��  ���F!�\a�} ��� ��� �� �� �� �� ��� ��� ��vz�MM�[�� ��  ��  ��  �����������������������������������d@@��  ��  ��  ��  �� �j�D3�Y]�ot�y }�| ��{ �w {�in�PP�G#���� ��  ��  ��  ��  �c??�������������������������������������a''��  ��  ��  ��  �� �� ���W�I$�F,�G*�L�a���� ��  ��  ��  ��  ��  �a&&���������������������������������������������d??����  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ���d>>���������������������������������������������������������hBB�p�~���������������������~�p�hAA����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
���
����                                                                                                                        ����(                                    ���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���������������������rr��qp��qo��qo��qp��rr����������������������������������!!��  ��  �� �� �� �� ��  ��  ��!!����������������������""��  ���qC�n k�t x�t w�mg�v9����  ��!!������������������  ���i\������ ��� ��� ��z ��kO����  ��������������ss��  �oG�| ���?���f��~ �� �� �� ��z ��x6��  ��rr����������qp�� �p p�~ ���Q������{ }�} �~ �� ��� ��lc�� ��po����������qo�� �w |�} ��P��֯���\���Z���,����� ��q t�� ��po����������qo�� �w |�} ��P��ױ���`���n��ԫ���2��~ ��q t�� ��po����������qp�� �p q�~ ���Q������y {�z |������b��~ ��md�� ��po����������ss��  �nI�{ ���N��ٵ���m���w��ԫ���1��y �x7��  ��rr��������������  ���i ]�����M���P���L���&��{��jQ����  ������������������  ��  ���oE�l k�r w�r v�l h�u<��	��  ��������������������������  ��  �� 	�� �� �� ��  ��  ������������������������������������nn��ml��mk��mk��ml��nn������������������������w���w���w���w���w���w���w���w���w���w���w���w���w���w���w���w��                                                          ��  